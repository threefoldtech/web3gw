module explorer

import freeflowuniverse.crystallib.rpcwebsocket { RpcWsClient }

pub struct Explorer {
	RpcWsClient
}