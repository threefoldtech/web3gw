module solution

pub enum Capacity {
	small
	medium
	large
	extra_large
}
