module tfgrid

import freeflowuniverse.crystallib.rpcwebsocket { RpcWsClient }

pub struct TFGridClient {
	RpcWsClient
}
