module main

import freeflowuniverse.crystallib.rpcwebsocket { RpcWsClient }

import threefoldtech.threebot.eth
import threefoldtech.threebot.explorer
import threefoldtech.threebot.stellar
import threefoldtech.threebot.tfchain
import threefoldtech.threebot.tfgrid
import threefoldtech.threebot.nostr
//ADD NEW CLIENTS HERE

import flag
import log
import os
import time

const (
	default_server_address = 'http://127.0.0.1:8080'
)


fn execute_rpcs(mut client RpcWsClient, mut logger log.Logger, mnemonic string) ! {
	// ADD YOUR CALLS HERE
}


fn main() {
	// This is some code that allows us to quickly create a commmand line tool with arguments. 
	mut fp := flag.new_flag_parser(os.args)
	fp.application('Welcome to the web3_proxy client. The web3_proxy client allows you to execute all remote procedure calls that the web3_proxy server can handle.')
	fp.limit_free_args(0, 0)!
	fp.description('')
	fp.skip_executable()
	mnemonic := fp.string('mnemonic', `m`, '', 'The mnemonic to be used to call any function')
	address := fp.string('address', `a`, '${default_server_address}', 'The address of the web3_proxy server to connect to.')
	debug_log := fp.bool('debug', 0, false, 'By setting this flag the client will print debug logs too.')
	_ := fp.finalize() or {
		eprintln(err)
		println(fp.usage())
		exit(1)
	}

	mut logger := log.Logger(&log.Log{
		level: if debug_log { .debug } else { .info }
	})

	mut myclient := rpcwebsocket.new_rpcwsclient(address, &logger) or {
		logger.error('Failed creating rpc websocket client: ${err}')
		exit(1)
	}
	_ := spawn myclient.run()
	execute_rpcs(mut myclient, mut logger, mnemonic) or {
		logger.error("Failed executing calls: $err")
		exit(1)
	}
}
