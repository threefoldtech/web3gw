module tfchain

pub struct {
	
}