module tfgrid

pub struct PresearchResult {
pub:
	name           string
	machine_ygg_ip string
	machine_ipv6   string
	machine_ipv4   string
}
