module solution

enum Capacity {
	small
	medium
	large
	extra_large
}
