module main

import freeflowuniverse.crystallib.rpcwebsocket { RpcWsClient }
import threefoldtech.threebot.nostr { CreateChannelInput, CreateChannelMessageInput, FetchChannelMessageInput }
import flag
import log
import os

const (
	default_server_address = 'ws://127.0.0.1:8080'
)

fn execute_rpcs(mut client RpcWsClient, mut logger log.Logger, secret string) ! {
	mut nostr_client := nostr.new(mut client)

	key := if secret == '' {
		k := nostr_client.generate_keypair()!
		logger.info('Key: ${k}')
		k
	} else {
		secret
	}

	nostr_client.load(key)!

	nostr_client.connect_to_relay('https://nostr01.grid.tf/')!

	channel_id := nostr_client.create_channel(CreateChannelInput{
		name: 'my chan'
		about: 'my about'
		picture: 'my pic'
	})!

	channels := nostr_client.list_channels()!
	logger.info('channels ${channels}')

	for i in 0 .. 10 {
		nostr_client.create_channel_message(CreateChannelMessageInput{
			content: 'my new message number ${i}'
			channel_id: channel_id
			message_id: 'some id'
			public_key: 'some pk'
		})!
	}

	messages := nostr_client.get_channel_message(FetchChannelMessageInput{
		channel_id: channel_id
	})!

	logger.info('channel messages: ${messages}')
}

fn main() {
	mut fp := flag.new_flag_parser(os.args)
	fp.application('Welcome to the web3_proxy client. The web3_proxy client allows you to execute all remote procedure calls that the web3_proxy server can handle.')
	fp.limit_free_args(0, 0)!
	fp.description('')
	fp.skip_executable()
	secret := fp.string('secret', `s`, '', 'The secret to use for nostr.')
	address := fp.string('address', `a`, '${default_server_address}', 'The address of the web3_proxy server to connect to.')
	debug_log := fp.bool('debug', 0, false, 'By setting this flag the client will print debug logs too.')
	_ := fp.finalize() or {
		eprintln(err)
		println(fp.usage())
		exit(1)
	}

	mut logger := log.Logger(&log.Log{
		level: if debug_log { .debug } else { .info }
	})

	mut myclient := rpcwebsocket.new_rpcwsclient(address, &logger) or {
		logger.error('Failed creating rpc websocket client: ${err}')
		exit(1)
	}

	_ := spawn myclient.run()

	execute_rpcs(mut myclient, mut logger, secret) or {
		logger.error('Failed executing calls: ${err}')
		exit(1)
	}
}
