module main

pub fn test(data string) int {
	println(data)
	return 0
}