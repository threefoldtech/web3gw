module zos

pub struct PublicIP4 {}

pub fn (p PublicIP4) challenge() string {
	return ''
}
