module threelang

// TFChainParser should handle all tfchain related actions
struct TFChainParser{

}