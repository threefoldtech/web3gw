module tfgrid

pub struct FunkwhaleResult {
pub:
	name           string
	machine_ygg_ip string
	machine_ipv6   string
	fqdn           string
}
