module tfgrid

pub struct TaigaResult {
pub:
	name           string
	machine_ygg_ip string
	machine_ipv6   string
	gateway_name   string
}
