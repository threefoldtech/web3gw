
module main

//TODO: import

import os

fn do()!{

//deploy 1 VM

}

fn main() {

	do() or {panic(err)}
}
