module threelang

// TFGridParser should handle parsing all tfgrid related actions
struct TFGridParser{

}